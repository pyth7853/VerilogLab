library verilog;
use verilog.vl_types.all;
entity FullAdd4 is
end FullAdd4;
